package ahb_package;
import uvm_pkg::*;
`include "uvm_macros.svh" 

  `include "ahb_sequence_item.sv"
  `include "ahb_sequence.sv"

  `include "ahb_driver.sv"
  `include "ahb_sequencer.sv"
  `include "ahb_agent.sv"
  `include "ahb_env.sv"


endpackage
